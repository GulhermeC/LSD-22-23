-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 17.1.0 Build 590 10/25/2017 SJ Lite Edition
-- Created on Tue May 09 15:00:24 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY DrinksFSM IS
    PORT (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        c : IN STD_LOGIC := '0';
        v : IN STD_LOGIC := '0';
        drink : OUT STD_LOGIC
    );
END DrinksFSM;

ARCHITECTURE BEHAVIOR OF DrinksFSM IS
    TYPE type_fstate IS (st0,st1,st2,st3,st4,st5);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clk,reg_fstate)
    BEGIN
        IF (clk='1' AND clk'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,c,v)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= st0;
            drink <= '0';
        ELSE
            drink <= '0';
            CASE fstate IS
                WHEN st0 =>
                    IF ((v = '1')) THEN
                        reg_fstate <= st1;
                    ELSIF ((NOT((v = '1')) AND (c = '1'))) THEN
                        reg_fstate <= st3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= st0;
                    END IF;

                    drink <= '0';
                WHEN st1 =>
                    IF ((v = '1')) THEN
                        reg_fstate <= st2;
                    ELSIF ((NOT((v = '1')) AND (c = '1'))) THEN
                        reg_fstate <= st4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= st1;
                    END IF;

                    drink <= '0';
                WHEN st2 =>
                    IF ((v = '1')) THEN
                        reg_fstate <= st3;
                    ELSIF ((NOT((v = '1')) AND (c = '1'))) THEN
                        reg_fstate <= st5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= st2;
                    END IF;

                    drink <= '0';
                WHEN st3 =>
                    IF ((v = '1')) THEN
                        reg_fstate <= st4;
                    ELSIF ((NOT((v = '1')) AND (c = '1'))) THEN
                        reg_fstate <= st5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= st3;
                    END IF;

                    drink <= '0';
                WHEN st4 =>
                    IF (((v = '1') OR (c = '1'))) THEN
                        reg_fstate <= st5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= st4;
                    END IF;

                    drink <= '0';
                WHEN st5 =>
                    reg_fstate <= st0;

                    drink <= '1';
                WHEN OTHERS => 
                    drink <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
