library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity DisplayDemoVHDL is
	port(	KEY 	: in std_logic_vector(0 downto 0);
			SW 	: in std_logic_vector (3 downto 0);
			HEX0	: out std_logic_vector (6 downto 0);
			LEDG	: out std_logic_vector (3 downto 0);
			LEDR	: out std_logic_vector (6 downto 0));
end DisplayDemoVHDL;

architecture Shell of DisplayDemoVHDL is
signal s_aulixiar : std_logic_vector(6 downto 0);

begin
	Disp : entity work.Bin7SegDecoder(Behavioral)
					port map(enable 	=> KEY(0),
								binInput => SW,
								decOut_n => s_aulixiar);
	
	HEX0(6 downto 0) <= s_aulixiar;
	
	LEDG(3 downto 0) <= SW;
	
	LEDG(6 downto 0) <= s_aulixiar;
	

end Shell;